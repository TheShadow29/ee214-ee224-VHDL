--author :: Prof. Madhav Desai

entity lab5 is
   port(x1,x0,y1,y0: in bit;
        s1,s0: out bit);
end entity;

architecture Formulas of lab5 is
   signal w, z: bit;
begin
   s0 <= (y0 and (not x0)) or ((not y0) and x0);
   w  <= (y1 and (not x1)) or ((not y1) and x1);
   z  <= (y0 and x0);
   s1 <= (w  and (not z)) or ((not w) and z);
end Formulas;